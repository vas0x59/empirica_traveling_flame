THERMO
300.000   1000.000  5000.000

!000000
 GRI-Mech Version 3.0 Thermodynamics released 7/30/99
 NASA Polynomial format for CHEMKIN-II
 see README file for disclaimer
N2                      N   2               G300.000   5000.000  1000.000      1
 2.92664000E+00 1.48797680E-03-5.68476000E-07 1.00970380E-10-6.75335100E-15    2
-9.22797700E+02 5.98052800E+00 3.29867700E+00 1.40824040E-03-3.96322200E-06    3
 5.64151500E-09-2.44485400E-12-1.02089990E+03 3.95037200E+00                   4
AR                000000Ar  1               G300.000   5000.000  5000.000      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 4.36600000E+00 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 4.36600000E+00                   4
HE                000000He  1               G300.000   5000.000  5000.000      1
 2.50000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00 0.00000000E+00    2
-7.45375000E+02 9.28723974E-01 2.50000000E+00 0.00000000E+00 0.00000000E+00    3
 0.00000000E+00 0.00000000E+00-7.45375000E+02 9.28723974E-01                   4
H                 000000H   1               G300.000   5000.000  1000.000      1
 2.50000001E+00-2.30842973E-11 1.61561948E-14-4.73515235E-18 4.98197357E-22    2
 2.54736599E+04-4.46682914E-01 2.50000000E+00 7.05332819E-13-1.99591964E-15    3
 2.30081632E-18-9.27732332E-22 2.54736599E+04-4.46682853E-01                   4
O2                000000O   2               G300.000   5000.000  1000.000      1
 3.28253784E+00 1.48308754E-03-7.57966669E-07 2.09470555E-10-2.16717794E-14    2
-1.08845772E+03 5.45323129E+00 3.78245636E+00-2.99673416E-03 9.84730201E-06    3
-9.68129509E-09 3.24372837E-12-1.06394356E+03 3.65767573E+00                   4
OH                000000H   1O   1          G300.000   5000.000  1000.000      1
 2.86472886E+00 1.05650448E-03-2.59082758E-07 3.05218674E-11-1.33195876E-15    2
 3.71885774E+03 5.70164073E+00 4.12530561E+00-3.22544939E-03 6.52764691E-06    3
-5.79853643E-09 2.06237379E-12 3.38153812E+03-6.90432960E-01                   4
O                 000000O   1               G300.000   5000.000  1000.000      1
 2.56942078E+00-8.59741137E-05 4.19484589E-08-1.00177799E-11 1.22833691E-15    2
 2.92175791E+04 4.78433864E+00 3.16826710E+00-3.27931884E-03 6.64306396E-06    3
-6.12806624E-09 2.11265971E-12 2.91222592E+04 2.05193346E+00                   4
H2                000000H   2               G300.000   5000.000  1000.000      1
 3.33727920E+00-4.94024731E-05 4.99456778E-07-1.79566394E-10 2.00255376E-14    2
-9.50158922E+02-3.20502331E+00 2.34433112E+00 7.98052075E-03-1.94781510E-05    3
 2.01572094E-08-7.37611761E-12-9.17935173E+02 6.83010238E-01                   4
H2O               000000H   2O   1          G300.000   5000.000  1000.000      1
 3.03399249E+00 2.17691804E-03-1.64072518E-07-9.70419870E-11 1.68200992E-14    2
-3.00042971E+04 4.96677010E+00 4.19864056E+00-2.03643410E-03 6.52040211E-06    3
-5.48797062E-09 1.77197817E-12-3.02937267E+04-8.49032208E-01                   4
HO2               000000H   1O   2          G300.000   5000.000  1000.000      1
 4.01721090E+00 2.23982013E-03-6.33658150E-07 1.14246370E-10-1.07908535E-14    2
 1.11856713E+02 3.78510215E+00 4.30179801E+00-4.74912051E-03 2.11582891E-05    3
-2.42763894E-08 9.29225124E-12 2.94808040E+02 3.71666245E+00                   4
CO                000000C   1O   1          G300.000   5000.000  1000.000      1
 2.71518561E+00 2.06252743E-03-9.98825771E-07 2.30053008E-10-2.03647716E-14    2
-1.41518724E+04 7.81868772E+00 3.57953347E+00-6.10353680E-04 1.01681433E-06    3
 9.07005884E-10-9.04424499E-13-1.43440860E+04 3.50840928E+00                   4
CO2               000000C   1O   2          G300.000   5000.000  1000.000      1
 3.85746029E+00 4.41437026E-03-2.21481404E-06 5.23490188E-10-4.72084164E-14    2
-4.87591660E+04 2.27163806E+00 2.35677352E+00 8.98459677E-03-7.12356269E-06    3
 2.45919022E-09-1.43699548E-13-4.83719697E+04 9.90105222E+00                   4
HCO               000000C   1H   1O   1     G300.000   5000.000  1000.000      1
 2.77217438E+00 4.95695526E-03-2.48445613E-06 5.89161778E-10-5.33508711E-14    2
 4.01191815E+03 9.79834492E+00 4.22118584E+00-3.24392532E-03 1.37799446E-05    3
-1.33144093E-08 4.33768865E-12 3.83956496E+03 3.39437243E+00                   4
CH3               000000C   1H   3          G300.000   5000.000  1000.000      1
 2.28571772E+00 7.23990037E-03-2.98714348E-06 5.95684644E-10-4.67154394E-14    2
 1.67755843E+04 8.48007179E+00 3.67359040E+00 2.01095175E-03 5.73021856E-06    3
-6.87117425E-09 2.54385734E-12 1.64449988E+04 1.60456433E+00                   4
CH4               000000C   1H   4          G300.000   5000.000  1000.000      1
 7.48514950E-02 1.33909467E-02-5.73285809E-06 1.22292535E-09-1.01815230E-13    2
-9.46834459E+03 1.84373180E+01 5.14987613E+00-1.36709788E-02 4.91800599E-05    3
-4.84743026E-08 1.66693956E-11-1.02466476E+04-4.64130376E+00                   4
CH2O              000000C   1H   2O   1     G300.000   5000.000  1000.000      1
 1.76069008E+00 9.20000082E-03-4.42258813E-06 1.00641212E-09-8.83855640E-14    2
-1.39958323E+04 1.36563230E+01 4.79372315E+00-9.90833369E-03 3.73220008E-05    3
-3.79285261E-08 1.31772652E-11-1.43089567E+04 6.02812900E-01                   4
T-CH2             000000C   1H   2          G300.000   5000.000  1000.000      1
 2.87410113E+00 3.65639292E-03-1.40894597E-06 2.60179549E-10-1.87727567E-14    2
 4.62636040E+04 6.17119324E+00 3.76267867E+00 9.68872143E-04 2.79489841E-06    3
-3.85091153E-09 1.68741719E-12 4.60040401E+04 1.56253185E+00                   4
S-CH2             000000C   1H   2          G300.000   5000.000  1000.000      1
 2.29203842E+00 4.65588637E-03-2.01191947E-06 4.17906000E-10-3.39716365E-14    2
 5.09259997E+04 8.62650169E+00 4.19860411E+00-2.36661419E-03 8.23296220E-06    3
-6.68815981E-09 1.94314737E-12 5.04968163E+04-7.69118967E-01                   4
C2H4              000000C   2H   4          G300.000   5000.000  1000.000      1
 2.03611116E+00 1.46454151E-02-6.71077915E-06 1.47222923E-09-1.25706061E-13    2
 4.93988614E+03 1.03053693E+01 3.95920148E+00-7.57052247E-03 5.70990292E-05    3
-6.91588753E-08 2.69884373E-11 5.08977593E+03 4.09733096E+00                   4
CH3O              000000C   1H   3O   1     G300.000   5000.000  1000.000      1
 4.75779238E+00 7.44142474E-03-2.69705176E-06 4.38090504E-10-2.63537098E-14    2
 3.90139164E+02-1.96680028E+00 3.71180502E+00-2.80463306E-03 3.76550971E-05    3
-4.73072089E-08 1.86588420E-11 1.30772484E+03 6.57240864E+00                   4
C2H5              000000C   2H   5          G300.000   5000.000  1000.000      1
 1.95465642E+00 1.73972722E-02-7.98206668E-06 1.75217689E-09-1.49641576E-13    2
 1.28575200E+04 1.34624343E+01 4.30646568E+00-4.18658892E-03 4.97142807E-05    3
-5.99126606E-08 2.30509004E-11 1.28416265E+04 4.70720924E+00                   4
C2H6              000000C   2H   6          G300.000   5000.000  1000.000      1
 1.07188150E+00 2.16852677E-02-1.00256067E-05 2.21412001E-09-1.90002890E-13    2
-1.14263932E+04 1.51156107E+01 4.29142492E+00-5.50154270E-03 5.99438288E-05    3
-7.08466285E-08 2.68685771E-11-1.15222055E+04 2.66682316E+00                   4
H2O2              000000H   2O   2          G300.000   5000.000  1000.000      1
 4.16500285E+00 4.90831694E-03-1.90139225E-06 3.71185986E-10-2.87908305E-14    2
-1.78617877E+04 2.91615662E+00 4.27611269E+00-5.42822417E-04 1.67335701E-05    3
-2.15770813E-08 8.62454363E-12-1.77025821E+04 3.43505074E+00                   4
C2H2              000000C   2H   2          G300.000   5000.000  1000.000      1
 4.14756964E+00 5.96166664E-03-2.37294852E-06 4.67412171E-10-3.61235213E-14    2
 2.59359992E+04-1.23028121E+00 8.08681094E-01 2.33615629E-02-3.55171815E-05    3
 2.80152437E-08-8.50072974E-12 2.64289807E+04 1.39397051E+01                   4
C2H3              000000C   2H   3          G300.000   5000.000  1000.000      1
 3.01672400E+00 1.03302292E-02-4.68082349E-06 1.01763288E-09-8.62607041E-14    2
 3.46128739E+04 7.78732378E+00 3.21246645E+00 1.51479162E-03 2.59209412E-05    3
-3.57657847E-08 1.47150873E-11 3.48598468E+04 8.51054025E+00                   4
CH2CHO            000000C   2H   3O   1     G300.000   5000.000  1000.000      1
 5.16620060E+00 1.08478260E-02-4.46583680E-06 8.06285480E-10-4.84101930E-14    2
-7.31993470E+02-1.96333610E+00 1.01340010E+00 2.26814670E-02-1.57339440E-05    3
 4.04915030E-09 2.95990120E-13 3.80428530E+02 1.93565520E+01                   4
CH2CO             000000C   2H   2O   1     G300.000   5000.000  1000.000      1
 4.51129732E+00 9.00359745E-03-4.16939635E-06 9.23345882E-10-7.94838201E-14    2
-7.55105311E+03 6.32247205E-01 2.13583630E+00 1.81188721E-02-1.73947474E-05    3
 9.34397568E-09-2.01457615E-12-7.04291804E+03 1.22156480E+01                   4
CH2OH             000000C   1H   3O   1     G300.000   5000.000  1000.000      1
 5.09312037E+00 5.94758550E-03-2.06496524E-06 3.23006703E-10-1.88125052E-14    2
-4.05813228E+03-1.84690613E+00 4.47832317E+00-1.35069687E-03 2.78483707E-05    3
-3.64867397E-08 1.47906775E-11-3.52476728E+03 3.30911984E+00                   4
CH3CHO            000000C   2H   4O   1     G300.000   5000.000  1000.000      1
 5.40411080E+00 1.17230590E-02-4.22631370E-06 6.83724510E-10-4.09848630E-14    2
-2.25931220E+04-3.48079170E+00 4.72945950E+00-3.19328580E-03 4.75349210E-05    3
-5.74586110E-08 2.19311120E-11-2.15728780E+04 4.10301590E+00                   4
CH3CO             000000C   2H   3O   1     G300.000   5000.000  1000.000      1
 5.94477310E+00 7.86672050E-03-2.88658820E-06 4.72708750E-10-2.85998610E-14    2
-3.78730750E+03-5.01367510E+00 4.16342570E+00-2.32616100E-04 3.42678200E-05    3
-4.41052270E-08 1.72756120E-11-2.65745290E+03 7.34682800E+00                   4
C2H5OH            000000C   2H   6O   1     G300.000   5000.000  1000.000      1
 4.34717120E+00 1.86288000E-02-6.77946700E-06 8.16592600E-10 0.00000000E+00    2
-3.06615743E+04 3.24247304E+00 5.76535800E-01 2.89451200E-02-1.61002000E-05    3
 3.59164100E-09 0.00000000E+00-2.96359500E+04 2.27081300E+01                   4
CH2CH2OH          000000C   2H   5O   1     G300.000   5000.000  1000.000      1
 7.52244726E+00 1.10492715E-02-3.72576465E-06 5.72827397E-10-3.30061759E-14    2
-7.29337464E+03-1.24960750E+01 1.17714711E+00 2.48115685E-02-1.50299503E-05    3
 4.79006785E-09-6.40994211E-13-4.95369043E+03 2.20081586E+01                   4
CH3CHOH           000000C   2H   5O   1     G300.000   5000.000  1000.000      1
 7.26570301E+00 1.09588926E-02-3.63662803E-06 5.53659830E-10-3.17012322E-14    2
-8.64371441E+03-1.06822851E+01 1.83974631E+00 1.87789371E-02-4.60544253E-06    3
-2.13116990E-09 9.43772653E-13-6.29595195E+03 2.01446141E+01                   4
CH3CH2O           000000C   2H   5O   1     G300.000   5000.000  1000.000      1
 8.31182392E+00 1.03426319E-02-3.39186089E-06 5.12212617E-10-2.91601713E-14    2
-6.13097954E+03-2.13985581E+01-2.71296378E-01 2.98839812E-02-1.97090548E-05    3
 6.37339893E-09-7.77965054E-13-3.16397196E+03 2.47706003E+01                   4
END
